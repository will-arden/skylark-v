
module imem(
    
    input logic [31:0]      A,          // Address to read from
    output logic [31:0]     InstrF      // Output instruction
    
);

    

endmodule
