/*
Top-Level Module
-----------------
This module is the highest level in the project; all other modules are instantiated under here, including memories.
*/

module top_level();

rv_core rv_core;                // Instantiate the processor core

endmodule
